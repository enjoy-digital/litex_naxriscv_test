module NaxRiscvLitex (
  output              ram_ibus_arvalid,
  input               ram_ibus_arready,
  output     [31:0]   ram_ibus_araddr,
  output     [7:0]    ram_ibus_arlen,
  output     [2:0]    ram_ibus_arsize,
  output     [1:0]    ram_ibus_arburst,
  input               ram_ibus_rvalid,
  output              ram_ibus_rready,
  input      [63:0]   ram_ibus_rdata,
  input      [1:0]    ram_ibus_rresp,
  input               ram_ibus_rlast,
  output              ram_dbus_awvalid,
  input               ram_dbus_awready,
  output     [31:0]   ram_dbus_awaddr,
  output     [0:0]    ram_dbus_awid,
  output     [7:0]    ram_dbus_awlen,
  output     [2:0]    ram_dbus_awsize,
  output     [1:0]    ram_dbus_awburst,
  output              ram_dbus_wvalid,
  input               ram_dbus_wready,
  output     [63:0]   ram_dbus_wdata,
  output     [7:0]    ram_dbus_wstrb,
  output              ram_dbus_wlast,
  input               ram_dbus_bvalid,
  output              ram_dbus_bready,
  input      [0:0]    ram_dbus_bid,
  input      [1:0]    ram_dbus_bresp,
  output              ram_dbus_arvalid,
  input               ram_dbus_arready,
  output     [31:0]   ram_dbus_araddr,
  output     [0:0]    ram_dbus_arid,
  output     [7:0]    ram_dbus_arlen,
  output     [2:0]    ram_dbus_arsize,
  output     [1:0]    ram_dbus_arburst,
  input               ram_dbus_rvalid,
  output              ram_dbus_rready,
  input      [63:0]   ram_dbus_rdata,
  input      [0:0]    ram_dbus_rid,
  input      [1:0]    ram_dbus_rresp,
  input               ram_dbus_rlast,
  output              peripheral_ibus_arvalid,
  input               peripheral_ibus_arready,
  output     [31:0]   peripheral_ibus_araddr,
  output     [2:0]    peripheral_ibus_arprot,
  input               peripheral_ibus_rvalid,
  output              peripheral_ibus_rready,
  input      [63:0]   peripheral_ibus_rdata,
  input      [1:0]    peripheral_ibus_rresp,
  output              peripheral_dbus_awvalid,
  input               peripheral_dbus_awready,
  output     [31:0]   peripheral_dbus_awaddr,
  output     [2:0]    peripheral_dbus_awprot,
  output              peripheral_dbus_wvalid,
  input               peripheral_dbus_wready,
  output     [31:0]   peripheral_dbus_wdata,
  output     [3:0]    peripheral_dbus_wstrb,
  input               peripheral_dbus_bvalid,
  output              peripheral_dbus_bready,
  input      [1:0]    peripheral_dbus_bresp,
  output              peripheral_dbus_arvalid,
  input               peripheral_dbus_arready,
  output     [31:0]   peripheral_dbus_araddr,
  output     [2:0]    peripheral_dbus_arprot,
  input               peripheral_dbus_rvalid,
  output              peripheral_dbus_rready,
  input      [31:0]   peripheral_dbus_rdata,
  input      [1:0]    peripheral_dbus_rresp,
  input               peripheral_clint_CYC,
  input               peripheral_clint_STB,
  output              peripheral_clint_ACK,
  input               peripheral_clint_WE,
  input      [13:0]   peripheral_clint_ADR,
  output     [31:0]   peripheral_clint_DAT_MISO,
  input      [31:0]   peripheral_clint_DAT_MOSI,
  input               peripheral_plic_CYC,
  input               peripheral_plic_STB,
  output              peripheral_plic_ACK,
  input               peripheral_plic_WE,
  input      [21:0]   peripheral_plic_ADR,
  output     [31:0]   peripheral_plic_DAT_MISO,
  input      [31:0]   peripheral_plic_DAT_MOSI,
  input      [31:0]   peripheral_interrupt,
  input               clk,
  input               reset
);

endmodule